`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:27:55 02/05/2020 
// Design Name: 
// Module Name:    SR_FF 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SR_FF(S,R,clk,Q,Qbar
    );

input S,R,clk;
output reg Q,Qbar;

always@(posedge clk)
	begin
		Q<=S|((!R)&Q);
		Qbar<=R|((!S)&(!Q));
	end
endmodule
